// EASE/HDL begin //////////////////////////////////////////////////////////////
// 
// module 'LogicReset'.
// 
////////////////////////////////////////////////////////////////////////////////

module LogicReset (Rst, ReadyKey, RstKey) ;
  input      Rst;
  input      ReadyKey;
  output     RstKey;


// EASE/HDL end ////////////////////////////////////////////////////////////////



endmodule // LogicReset
